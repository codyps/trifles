.include "a1_fig.spice"

Vs  Vcc 0 DC 5v

*                PULSE(V1 V2 TD TR TF PW  PER)
Vi1 b_e1 0 DC 0  PULSE(0  5  0  2n 2n 0.5 1)
Vi0 a_e1 0 DC 0  PULSE(0  5  0  2n 2n 1   2)

.control

* .tran tstep tstop < tstart <tmax > > < uic >
tran 0.02 2
hardcopy a1_p1.eps v(a_e1) v(b_e1) v(c3) 


.endc
.enc
