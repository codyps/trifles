* Lab 2, Act 1, NMOS inverter, #6

.include 'nmos_inv_broken.spice'

nmos_inv 0 vin_r vout vdd

rin vin vin_r 1k
Vsdd vdd 0 DC 5
Vsin vin 0 DC 0

.control
dc Vsin 0 5 0.01
hardcopy p1.eps V(vout) V(vin)
.endc
.end
