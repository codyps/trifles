`include "p11_12.v"

module a16_test();
	/* as we can assume that the 4bit adder was succesfully tested, our
	 * goal here is simply to cause the carry interconects (of which there
	 * are 4) to triger in all possible arrangments (16)
	 */

	reg ra1[3:0], ra2[3:0], ra3[3:0], ra4[3:0];
	reg rb1[3:0], rb2[3:0], rb3[3:0], rb4[3:0];


	initial begin


	end
endmodule
