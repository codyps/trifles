* a4_p1.spice
.include 'a3_fig.spice'

Vs  Vee  0 -1.8
Vsr Vref 0 -1.2

*                PULSE(V1 V2 TD TR TF PW  PER)
Vi0 0 A PULSE(0  1.6  0  2n 2n 0.5 1)
Vi1 0 B PULSE(0  1.6  0  2n 2n 1   2)

.control

* .tran tstep tstop < tstart <tmax > > < uic >
tran 0.02 2
hardcopy include/a4_p1.eps v(A) v(B) v(OR) 

.endc
.end
