* a4_p2.spice
.include "a3_fig.spice"

Vs  0 Vee  DC 1.8
Vsr 0 Vref DC 1.2

Vi0 0 A DC 1.6
Vi1 0 B

.control
* .dc srcnam vstart vstop vincr [ src2 start2 stop2 incr2 ]
dc Vi1 0.8 1.8 0.1
hardcopy include/a4_p2.eps v(B) v(OR) 
.endc
.end
