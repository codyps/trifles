.include "Q2N3904.spice"
.include "DN4001.spice"

RB1 Vcc b1 4k
RB2 Vcc b2 4k

RC1 Vcc c3 1.5k
RC2 Vcc c6 120

RE  e4 0 1k

*  C  B  E
Q1 c1 b1 A  Q2N3904
Q2 c2 b2 B  Q2N3904
Q3 c3 c1 e3 Q2N3904
Q4 c4 c2 e3 Q2N3904
Q5 Y  e3 0  Q2N3904

D1 0 A DN4001
D2 0 B DN4001

