
.MODEL  DN4001  D  (IS=5.86E-06 N=1.7 BV=6.66E+1 IBV=5.0E-07
+ RS=3.62E-02 CJO=5.21E-11 VJ=.34 M=.38 TT=5.04E-06)
