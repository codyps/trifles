* Normal nmos inverter.

.subckt nmos_inv gnd vin vout vdd
Ml  vdd  vdd vout gnd NMOS
Msa vout vin gnd  gnd NMOS
Msb vout vin gnd  gnd NMOS
.ends
