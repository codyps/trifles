.include "a2_fig.spice"

Vs  Vcc 0 DC 5v

*                PULSE(V1 V2 TD TR TF PW  PER)
Vi0 A 0 DC 0  PULSE(0  5  0  2n 2n 0.5 1)
Vi1 B 0 DC 0  PULSE(0  5  0  2n 2n 1   2)

.control

* .tran tstep tstop < tstart <tmax > > < uic >
tran 0.02 2
hardcopy include/a2_p1.eps v(A) v(B) v(Y) 

.endc
.enc
