module Y1(output Y, input A,B,C,D);
	//Σm (4,5,6,7,11,12,13)
	
endmodule

module Y2(output Y, input A,B,C,D);
	//Σm (1,2,3,4)
endmodule
