
* .model IRF150
* + NMOS(Level=3 Gamma=0 Delta=0 Eta=0 Theta=0 Kappa=0 Vmax=0 Xj=0
* +Tox=100n Uo=600 Phi=.6 Rs=1.624m Kp=50u W=160u L=2u Vto=2
* +Rd=1.031m Rds=444.4K Cbd=3.229n Pb=.8 Mj=.5 Fc=.5 Cgso=9.027n
* +Cgdo=1.679n Rg=13.89 Is=194E-18 N=1 Tt=288n lambda=0.05)
* * Int'l Rectifier pid=IRFC150 case=TO3 88-08-25 bam creation

.model irf150 nmos (TOX=100N PHI=.6 KP=20.53U W=.3
+ L=2U VTO=2.831 RD=1.031M RDS=444.4K CBD=3.229N
+ PB=.8 MJ=.5
+ CGSO=9.027N CGDO=1.679N RG=13.89 IS=194e-18 N=1
+ TT=288N)



