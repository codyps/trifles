.include "Q2N3904.spice"

RC1 0 b4 270
RC2 0 b3 300

RE1 ea  Vee 1.2k
RE2 OR  Vee 2k
RE3 NOR Vee 2k

*   C  B    E
Q1A b4 A    ea
Q1B b4 B    ea
Q2  b3 Vref ea
Q3  0  b3   OR
Q4  0  b4   NOR
